magic
tech sky130A
magscale 1 2
timestamp 1652441850
<< nwell >>
rect 309 466 731 1234
<< pwell >>
rect 309 -95 731 463
<< nmos >>
rect 505 53 535 253
<< pmos >>
rect 505 686 535 1086
<< ndiff >>
rect 447 241 505 253
rect 447 65 459 241
rect 493 65 505 241
rect 447 53 505 65
rect 535 241 593 253
rect 535 65 547 241
rect 581 65 593 241
rect 535 53 593 65
<< pdiff >>
rect 447 1074 505 1086
rect 447 698 459 1074
rect 493 698 505 1074
rect 447 686 505 698
rect 535 1074 593 1086
rect 535 698 547 1074
rect 581 698 593 1074
rect 535 686 593 698
<< ndiffc >>
rect 459 65 493 241
rect 547 65 581 241
<< pdiffc >>
rect 459 698 493 1074
rect 547 698 581 1074
<< psubdiff >>
rect 345 393 441 427
rect 599 393 695 427
rect 345 331 379 393
rect 661 331 695 393
rect 345 -25 379 37
rect 661 -25 695 37
rect 345 -59 441 -25
rect 599 -59 695 -25
<< nsubdiff >>
rect 345 1164 441 1198
rect 599 1164 695 1198
rect 345 1101 379 1164
rect 661 1101 695 1164
rect 345 536 379 599
rect 661 536 695 599
rect 345 502 441 536
rect 599 502 695 536
<< psubdiffcont >>
rect 441 393 599 427
rect 345 37 379 331
rect 661 37 695 331
rect 441 -59 599 -25
<< nsubdiffcont >>
rect 441 1164 599 1198
rect 345 599 379 1101
rect 661 599 695 1101
rect 441 502 599 536
<< poly >>
rect 505 1086 535 1112
rect 505 655 535 686
rect 487 639 553 655
rect 487 605 503 639
rect 537 605 553 639
rect 487 589 553 605
rect 487 325 553 341
rect 487 291 503 325
rect 537 291 553 325
rect 487 275 553 291
rect 505 253 535 275
rect 505 27 535 53
<< polycont >>
rect 503 605 537 639
rect 503 291 537 325
<< locali >>
rect 345 1164 441 1198
rect 599 1164 695 1198
rect 345 1101 379 1164
rect 661 1101 695 1164
rect 459 1074 493 1090
rect 459 682 493 698
rect 547 1074 581 1090
rect 547 682 581 698
rect 487 605 503 639
rect 537 605 553 639
rect 345 536 379 599
rect 661 536 695 599
rect 345 502 441 536
rect 599 502 695 536
rect 345 393 441 427
rect 599 393 695 427
rect 345 331 379 393
rect 661 331 695 393
rect 487 291 503 325
rect 537 291 553 325
rect 459 241 493 257
rect 459 49 493 65
rect 547 241 581 257
rect 547 49 581 65
rect 345 -25 379 37
rect 661 -25 695 37
rect 345 -59 441 -25
rect 599 -59 695 -25
<< viali >>
rect 345 826 379 957
rect 459 698 493 1074
rect 547 698 581 1074
rect 503 605 537 639
rect 503 291 537 325
rect 345 117 379 205
rect 459 65 493 241
rect 547 65 581 241
<< metal1 >>
rect 453 1074 499 1086
rect 51 903 251 991
rect 339 957 385 969
rect 339 903 345 957
rect 51 871 345 903
rect 51 791 251 871
rect 339 826 345 871
rect 379 903 385 957
rect 453 903 459 1074
rect 379 871 459 903
rect 379 826 385 871
rect 339 814 385 826
rect 453 698 459 871
rect 493 698 499 1074
rect 453 686 499 698
rect 541 1074 587 1086
rect 541 698 547 1074
rect 581 906 587 1074
rect 581 861 737 906
rect 581 698 587 861
rect 541 686 587 698
rect 491 639 549 645
rect 491 605 503 639
rect 537 605 549 639
rect 63 483 263 570
rect 491 483 549 605
rect 63 449 549 483
rect 63 370 263 449
rect 491 325 549 449
rect 491 291 503 325
rect 537 291 549 325
rect 491 285 549 291
rect 703 481 737 861
rect 767 481 967 573
rect 703 450 967 481
rect 453 241 499 253
rect 159 181 270 215
rect 339 205 385 217
rect 339 181 345 205
rect 159 141 345 181
rect 159 104 270 141
rect 339 117 345 141
rect 379 181 385 205
rect 453 181 459 241
rect 379 141 459 181
rect 379 117 385 141
rect 339 105 385 117
rect 453 65 459 141
rect 493 65 499 241
rect 453 53 499 65
rect 541 241 587 253
rect 541 65 547 241
rect 581 179 587 241
rect 703 179 737 450
rect 767 373 967 450
rect 581 134 737 179
rect 581 65 587 134
rect 703 133 737 134
rect 541 53 587 65
<< labels >>
flabel metal1 51 791 251 991 0 FreeSans 256 0 0 0 VDD
port 2 nsew
flabel metal1 63 370 263 570 0 FreeSans 256 0 0 0 A
port 0 nsew
flabel metal1 767 373 967 573 0 FreeSans 256 0 0 0 Y
port 1 nsew
flabel metal1 166 113 263 202 1 FreeSerif 160 0 0 0 VSS
port 3 n
<< end >>
